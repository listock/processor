/** CU testing suit.
 *
 * Author: Aleksandr Novozhilov
 * Creating date: 2018-06-14
 */

`include "cu.sv"

module cu_tb();

        initial begin
                $display("[CONTROL UNIT] test suit starts...");
                $display("[CONTROL UNIT] test suit ends.");
        end

endmodule